`timescale 1ns / 1ps

// This module forwards information
module Forward();
endmodule
